	"pnpm": {
		"onlyBuiltDependencies": [
		// 	"better-sqlite3",
		// 	"esbuild"
		 ]
	},
